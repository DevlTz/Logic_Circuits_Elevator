-- ean, não fiz ainda, mas vamo fzr depois! :)